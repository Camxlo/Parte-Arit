LIBRARY ieee;
USE ieee.std_logic_1164.all; 

LIBRARY work;

ENTITY Mux_Cuadru IS 
	PORT
	(
		A0 :  IN  STD_LOGIC;
		B0 :  IN  STD_LOGIC;
		A1 :  IN  STD_LOGIC;
		B1 :  IN  STD_LOGIC;
		A2 :  IN  STD_LOGIC;
		B2 :  IN  STD_LOGIC;
		A3 :  IN  STD_LOGIC;
		B3 :  IN  STD_LOGIC;
		S0 :  IN  STD_LOGIC;
		Y0 :  OUT  STD_LOGIC;
		Y1 :  OUT  STD_LOGIC;
		Y2 :  OUT  STD_LOGIC;
		Y3 :  OUT  STD_LOGIC
	);
END Mux_Cuadru;

ARCHITECTURE Part_Arit OF Mux_Cuadru IS 

SIGNAL	SYNTHESIZED_WIRE_0 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_1 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_17 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_3 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_4 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_6 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_7 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_18 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_15 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_16 :  STD_LOGIC;


BEGIN 



Y0 <= SYNTHESIZED_WIRE_0 OR SYNTHESIZED_WIRE_1;


SYNTHESIZED_WIRE_18 <= NOT(SYNTHESIZED_WIRE_17);



Y1 <= SYNTHESIZED_WIRE_3 OR SYNTHESIZED_WIRE_4;


SYNTHESIZED_WIRE_7 <= A0 AND SYNTHESIZED_WIRE_17;


Y3 <= SYNTHESIZED_WIRE_6 OR SYNTHESIZED_WIRE_7;


SYNTHESIZED_WIRE_6 <= B0 AND SYNTHESIZED_WIRE_18;


SYNTHESIZED_WIRE_16 <= A1 AND SYNTHESIZED_WIRE_17;


SYNTHESIZED_WIRE_15 <= B1 AND SYNTHESIZED_WIRE_18;


SYNTHESIZED_WIRE_4 <= A2 AND SYNTHESIZED_WIRE_17;


SYNTHESIZED_WIRE_3 <= B2 AND SYNTHESIZED_WIRE_18;


SYNTHESIZED_WIRE_1 <= A3 AND SYNTHESIZED_WIRE_17;


SYNTHESIZED_WIRE_0 <= B3 AND SYNTHESIZED_WIRE_18;


SYNTHESIZED_WIRE_17 <= NOT(S0);



Y2 <= SYNTHESIZED_WIRE_15 OR SYNTHESIZED_WIRE_16;


END Part_Arit;