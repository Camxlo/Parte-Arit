LIBRARY ieee;
USE ieee.std_logic_1164.all; 

LIBRARY work;

ENTITY FA IS 
	PORT
	(
		A :  IN  STD_LOGIC;
		B :  IN  STD_LOGIC;
		Cin :  IN  STD_LOGIC;
		Suma :  OUT  STD_LOGIC;
		Carry :  OUT  STD_LOGIC
	);
END FA;

ARCHITECTURE Part_Arit OF FA IS 

SIGNAL	SYNTHESIZED_WIRE_0 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_1 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_2 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_3 :  STD_LOGIC;


BEGIN 



SYNTHESIZED_WIRE_0 <= A XOR B;


Suma <= SYNTHESIZED_WIRE_0 XOR Cin;


SYNTHESIZED_WIRE_3 <= A AND B;


SYNTHESIZED_WIRE_1 <= B AND Cin;


SYNTHESIZED_WIRE_2 <= A AND Cin;


Carry <= SYNTHESIZED_WIRE_1 OR SYNTHESIZED_WIRE_2 OR SYNTHESIZED_WIRE_3;


END Part_Arit;